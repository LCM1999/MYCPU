library verilog;
use verilog.vl_types.all;
entity MyCPU is
    port(
        CLK             : in     vl_logic;
        RST             : in     vl_logic;
        nextPC          : out    vl_logic_vector(31 downto 0);
        currPC          : out    vl_logic_vector(31 downto 0);
        InsData         : out    vl_logic_vector(31 downto 0);
        IRIns           : out    vl_logic_vector(31 downto 0);
        op              : out    vl_logic_vector(5 downto 0);
        rs              : out    vl_logic_vector(4 downto 0);
        rt              : out    vl_logic_vector(4 downto 0);
        rd              : out    vl_logic_vector(4 downto 0);
        ID_immediate    : out    vl_logic_vector(15 downto 0);
        RegWre          : out    vl_logic;
        RegDst          : out    vl_logic;
        J               : out    vl_logic_vector(1 downto 0);
        MEM_Read        : out    vl_logic;
        MEM_Write       : out    vl_logic;
        MEMtoReg        : out    vl_logic;
        ExtSign         : out    vl_logic;
        ALUOp           : out    vl_logic_vector(2 downto 0);
        Reg_DataBusA    : out    vl_logic_vector(31 downto 0);
        Reg_DataBusB    : out    vl_logic_vector(31 downto 0);
        addr            : out    vl_logic_vector(4 downto 0);
        extended        : out    vl_logic_vector(31 downto 0);
        MEM_Con         : out    vl_logic_vector(1 downto 0);
        WB_Con          : out    vl_logic_vector(1 downto 0);
        ALUCon          : out    vl_logic_vector(2 downto 0);
        ID_EX_Reg_RS    : out    vl_logic_vector(4 downto 0);
        ID_EX_Reg_RT    : out    vl_logic_vector(4 downto 0);
        ID_EX_Reg_RD    : out    vl_logic_vector(4 downto 0);
        ID_EX_Reg_immediate: out    vl_logic_vector(31 downto 0);
        ID_EX_DataBusA  : out    vl_logic_vector(31 downto 0);
        ID_EX_DataBusB  : out    vl_logic_vector(31 downto 0);
        result          : out    vl_logic_vector(31 downto 0);
        EX_MEM_Write_Con: out    vl_logic;
        EX_MEM_Read_Con : out    vl_logic;
        EX_MEM_ALUOut   : out    vl_logic_vector(31 downto 0);
        EX_MEM_MEMtoReg : out    vl_logic;
        EX_MEM_RegWre   : out    vl_logic;
        EX_MEM_Reg_RD   : out    vl_logic_vector(4 downto 0);
        rData           : out    vl_logic_vector(31 downto 0);
        WB_RegWre       : out    vl_logic;
        WB_DataBus      : out    vl_logic_vector(31 downto 0);
        WB_Reg_RD       : out    vl_logic_vector(4 downto 0);
        stall           : out    vl_logic;
        ForwardA        : out    vl_logic_vector(1 downto 0);
        ForwardB        : out    vl_logic_vector(1 downto 0);
        Flash           : out    vl_logic;
        PCSrc           : out    vl_logic_vector(1 downto 0)
    );
end MyCPU;
