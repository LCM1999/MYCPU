library verilog;
use verilog.vl_types.all;
entity TestMyCPU is
end TestMyCPU;
